eefrf
