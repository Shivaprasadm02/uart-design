fde3frfg
