rfr43gf
